module ALU( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [3:0]  io_ALUOp, // @[:@6.4]
  input  [63:0] io_inputA, // @[:@6.4]
  input  [63:0] io_inputB, // @[:@6.4]
  output [63:0] io_output // @[:@6.4]
);
  wire [5:0] shamt; // @[alu.scala 27:26:@8.4]
  wire [64:0] _T_19; // @[alu.scala 35:37:@9.4]
  wire [63:0] _T_20; // @[alu.scala 35:37:@10.4]
  wire [63:0] _T_22; // @[alu.scala 36:37:@11.4]
  wire [63:0] _T_24; // @[alu.scala 37:37:@12.4]
  wire [63:0] _T_26; // @[alu.scala 38:37:@13.4]
  wire  _T_28; // @[alu.scala 39:38:@14.4]
  wire [126:0] _GEN_0; // @[alu.scala 40:37:@15.4]
  wire [126:0] _T_30; // @[alu.scala 40:37:@15.4]
  wire [63:0] _T_32; // @[alu.scala 41:37:@16.4]
  wire [63:0] _T_34; // @[alu.scala 42:38:@17.4]
  wire [63:0] _T_35; // @[alu.scala 42:45:@18.4]
  wire [63:0] _T_36; // @[alu.scala 42:55:@19.4]
  wire  _T_37; // @[Mux.scala 46:19:@20.4]
  wire [63:0] _T_38; // @[Mux.scala 46:16:@21.4]
  wire  _T_39; // @[Mux.scala 46:19:@22.4]
  wire [63:0] _T_40; // @[Mux.scala 46:16:@23.4]
  wire  _T_41; // @[Mux.scala 46:19:@24.4]
  wire [126:0] _T_42; // @[Mux.scala 46:16:@25.4]
  wire  _T_43; // @[Mux.scala 46:19:@26.4]
  wire [126:0] _T_44; // @[Mux.scala 46:16:@27.4]
  wire  _T_45; // @[Mux.scala 46:19:@28.4]
  wire [126:0] _T_46; // @[Mux.scala 46:16:@29.4]
  wire  _T_47; // @[Mux.scala 46:19:@30.4]
  wire [126:0] _T_48; // @[Mux.scala 46:16:@31.4]
  wire  _T_49; // @[Mux.scala 46:19:@32.4]
  wire [126:0] _T_50; // @[Mux.scala 46:16:@33.4]
  wire  _T_51; // @[Mux.scala 46:19:@34.4]
  wire [126:0] _T_52; // @[Mux.scala 46:16:@35.4]
  wire  _T_53; // @[Mux.scala 46:19:@36.4]
  wire [126:0] _T_54; // @[Mux.scala 46:16:@37.4]
  wire  _T_55; // @[Mux.scala 46:19:@38.4]
  wire [126:0] _T_56; // @[Mux.scala 46:16:@39.4]
  wire  _T_57; // @[Mux.scala 46:19:@40.4]
  wire [126:0] _T_58; // @[Mux.scala 46:16:@41.4]
  assign shamt = io_inputB[5:0]; // @[alu.scala 27:26:@8.4]
  assign _T_19 = io_inputA + io_inputB; // @[alu.scala 35:37:@9.4]
  assign _T_20 = io_inputA + io_inputB; // @[alu.scala 35:37:@10.4]
  assign _T_22 = io_inputA & io_inputB; // @[alu.scala 36:37:@11.4]
  assign _T_24 = io_inputA | io_inputB; // @[alu.scala 37:37:@12.4]
  assign _T_26 = io_inputA ^ io_inputB; // @[alu.scala 38:37:@13.4]
  assign _T_28 = io_inputA < io_inputB; // @[alu.scala 39:38:@14.4]
  assign _GEN_0 = {{63'd0}, io_inputA}; // @[alu.scala 40:37:@15.4]
  assign _T_30 = _GEN_0 << shamt; // @[alu.scala 40:37:@15.4]
  assign _T_32 = io_inputA >> shamt; // @[alu.scala 41:37:@16.4]
  assign _T_34 = $signed(io_inputA); // @[alu.scala 42:38:@17.4]
  assign _T_35 = $signed(_T_34) >>> shamt; // @[alu.scala 42:45:@18.4]
  assign _T_36 = $unsigned(_T_35); // @[alu.scala 42:55:@19.4]
  assign _T_37 = 4'ha == io_ALUOp; // @[Mux.scala 46:19:@20.4]
  assign _T_38 = _T_37 ? _T_36 : 64'h0; // @[Mux.scala 46:16:@21.4]
  assign _T_39 = 4'h9 == io_ALUOp; // @[Mux.scala 46:19:@22.4]
  assign _T_40 = _T_39 ? _T_32 : _T_38; // @[Mux.scala 46:16:@23.4]
  assign _T_41 = 4'h8 == io_ALUOp; // @[Mux.scala 46:19:@24.4]
  assign _T_42 = _T_41 ? _T_30 : {{63'd0}, _T_40}; // @[Mux.scala 46:16:@25.4]
  assign _T_43 = 4'h7 == io_ALUOp; // @[Mux.scala 46:19:@26.4]
  assign _T_44 = _T_43 ? {{126'd0}, _T_28} : _T_42; // @[Mux.scala 46:16:@27.4]
  assign _T_45 = 4'h6 == io_ALUOp; // @[Mux.scala 46:19:@28.4]
  assign _T_46 = _T_45 ? {{63'd0}, _T_26} : _T_44; // @[Mux.scala 46:16:@29.4]
  assign _T_47 = 4'h5 == io_ALUOp; // @[Mux.scala 46:19:@30.4]
  assign _T_48 = _T_47 ? {{63'd0}, _T_24} : _T_46; // @[Mux.scala 46:16:@31.4]
  assign _T_49 = 4'h4 == io_ALUOp; // @[Mux.scala 46:19:@32.4]
  assign _T_50 = _T_49 ? {{63'd0}, _T_22} : _T_48; // @[Mux.scala 46:16:@33.4]
  assign _T_51 = 4'h3 == io_ALUOp; // @[Mux.scala 46:19:@34.4]
  assign _T_52 = _T_51 ? {{63'd0}, _T_20} : _T_50; // @[Mux.scala 46:16:@35.4]
  assign _T_53 = 4'h2 == io_ALUOp; // @[Mux.scala 46:19:@36.4]
  assign _T_54 = _T_53 ? {{63'd0}, io_inputB} : _T_52; // @[Mux.scala 46:16:@37.4]
  assign _T_55 = 4'h1 == io_ALUOp; // @[Mux.scala 46:19:@38.4]
  assign _T_56 = _T_55 ? {{63'd0}, io_inputA} : _T_54; // @[Mux.scala 46:16:@39.4]
  assign _T_57 = 4'h0 == io_ALUOp; // @[Mux.scala 46:19:@40.4]
  assign _T_58 = _T_57 ? 127'h0 : _T_56; // @[Mux.scala 46:16:@41.4]
  assign io_output = _T_58[63:0]; // @[alu.scala 28:15:@42.4]
endmodule
